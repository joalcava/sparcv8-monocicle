----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    16:24:13 10/06/2016 
-- Design Name: 
-- Module Name:    Sparcv8Monocicle - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity Sparcv8Monocicle is
end Sparcv8Monocicle;

architecture Behavioral of Sparcv8Monocicle is

begin


end Behavioral;

