library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity sign_ext_unit is
end sign_ext_unit;

architecture Behavioral of sign_ext_unit is

begin


end Behavioral;

